///////////////////////////////////////////////////////////////////////////////////////////////////
//
// UVM SPI MEM TB pkg
// 
// This is the top level SPIMEM testbench package 
// SPI MEM
//
///////////////////////////////////////////////////////////////////////////////////////////////////

 package spi_mem_tb_pkg;
 
  import uvm_spi_mem_tests_pkg::*;
  
 endpackage